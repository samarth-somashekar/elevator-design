��` t i m e s c a l e   1 n s   /   1 p s  
  
 m o d u l e   E l e v a t o r 2 (  
         i n p u t   l o g i c   c l k ,   r e s e t ,  
         i n p u t   l o g i c   [ 4 : 0 ]   f l o o r _ r e q u e s t ,  
         o u t p u t   l o g i c   [ 4 : 0 ]   c u r r e n t _ f l o o r ,  
         o u t p u t   l o g i c   m o v i n g ,   d i r e c t i o n  
 ) ;  
  
         l o g i c   [ 2 : 0 ]   f r ,   c f ;  
         l o g i c   v a l i d _ r e q u e s t ;  
          
         l o g i c   c l k b i t ;  
         l o g i c   [ 2 7 : 0 ] c o u n t ;  
         a l w a y s _ f f @ ( p o s e d g e   c l k )  
         b e g i n  
                 c o u n t   < =   c o u n t   +   1 ;  
                 c l k b i t   =   c o u n t [ 2 7 ] ;  
         e n d  
          
         p r i o r i t y _ e n c o d e r   p r e ( . i p e ( f l o o r _ r e q u e s t ) ,   . o p e ( f r ) ,   . v a l i d ( v a l i d _ r e q u e s t ) ) ;  
  
         d e c o d e r   d e c ( . i p d ( c f ) ,   . o p d ( c u r r e n t _ f l o o r ) ) ;  
  
         a l w a y s _ f f   @ ( p o s e d g e   c o u n t [ 2 7 ]   o r   p o s e d g e   r e s e t )   b e g i n  
                 i f   ( r e s e t )   b e g i n  
                         c f   < =   3 ' d 0 ;  
                         m o v i n g   < =   0 ;  
                         d i r e c t i o n   < =   1 ;  
                 e n d    
                 e l s e   i f   ( v a l i d _ r e q u e s t )   b e g i n      
                         i f   ( c f   = =   f r )   b e g i n  
                                 m o v i n g   < =   0 ;            
                         e n d    
                         e l s e   b e g i n  
                                 m o v i n g   < =   1 ;            
                                 i f   ( c f   <   f r )   b e g i n  
                                         d i r e c t i o n   < =   1 ;      
                                         c f   < =   c f   +   1 ;  
                                 e n d    
                                 e l s e   b e g i n  
                                         d i r e c t i o n   < =   0 ;      
                                         c f   < =   c f   -   1 ;  
                                 e n d  
                         e n d  
                 e n d    
                 e l s e    
                         m o v i n g   < =   0 ;  
         e n d  
 e n d m o d u l e  
  
 m o d u l e   p r i o r i t y _ e n c o d e r (  
         i n p u t   l o g i c   [ 4 : 0 ]   i p e ,  
         o u t p u t   l o g i c   [ 2 : 0 ]   o p e ,  
         o u t p u t   l o g i c   v a l i d  
 ) ;  
         a l w a y s _ c o m b   b e g i n  
                 c a s e x   ( i p e )  
                         5 ' b 0 0 0 0 1   :   b e g i n   o p e   =   3 ' b 0 0 0 ;   v a l i d   =   1 ;   e n d  
                         5 ' b 0 0 0 1 x   :   b e g i n   o p e   =   3 ' b 0 0 1 ;   v a l i d   =   1 ;   e n d  
                         5 ' b 0 0 1 x x   :   b e g i n   o p e   =   3 ' b 0 1 0 ;   v a l i d   =   1 ;   e n d  
                         5 ' b 0 1 x x x   :   b e g i n   o p e   =   3 ' b 0 1 1 ;   v a l i d   =   1 ;   e n d  
                         5 ' b 1 x x x x   :   b e g i n   o p e   =   3 ' b 1 0 0 ;   v a l i d   =   1 ;   e n d  
                         d e f a u l t     :   b e g i n   o p e   =   3 ' b 0 0 0 ;   v a l i d   =   0 ;   e n d    
                 e n d c a s e  
         e n d  
 e n d m o d u l e  
  
 m o d u l e   d e c o d e r (  
         i n p u t   l o g i c   [ 2 : 0 ]   i p d ,  
         o u t p u t   l o g i c   [ 4 : 0 ]   o p d  
 ) ;  
         a l w a y s _ c o m b   b e g i n  
                 c a s e   ( i p d )  
                         3 ' b 0 0 0   :   o p d   =   5 ' b 0 0 0 0 1 ;  
                         3 ' b 0 0 1   :   o p d   =   5 ' b 0 0 0 1 0 ;  
                         3 ' b 0 1 0   :   o p d   =   5 ' b 0 0 1 0 0 ;  
                         3 ' b 0 1 1   :   o p d   =   5 ' b 0 1 0 0 0 ;  
                         3 ' b 1 0 0   :   o p d   =   5 ' b 1 0 0 0 0 ;  
                         d e f a u l t :   o p d   =   5 ' b 0 0 0 0 0 ;  
                 e n d c a s e  
         e n d  
 e n d m o d u l e  
 