�� 
 ` t i m e s c a l e   1 n s   /   1 p s  
  
 m o d u l e   E l e v a t o r 2 _ T B ( ) ;  
         l o g i c   c l k ,   r e s e t ;  
         l o g i c   [ 4 : 0 ]   f l o o r _ r e q u e s t ;  
         l o g i c   [ 4 : 0 ]   c u r r e n t _ f l o o r ;  
         l o g i c   m o v i n g ,   d i r e c t i o n ;  
          
         E l e v a t o r 2   d u t ( . c l k ( c l k ) ,   . r e s e t ( r e s e t ) ,   . f l o o r _ r e q u e s t ( f l o o r _ r e q u e s t ) ,   . c u r r e n t _ f l o o r ( c u r r e n t _ f l o o r ) ,   . m o v i n g ( m o v i n g ) ,   . d i r e c t i o n ( d i r e c t i o n ) ) ;  
          
         i n i t i a l    
         b e g i n  
                 f o r e v e r   # 5   c l k   =   ~ c l k ;  
         e n d  
          
         i n i t i a l    
         b e g i n  
         c l k   =   0 ;  
                 r e s e t   =   1 ;  
                 f l o o r _ r e q u e s t   =   5 ' b 1 0 0 0 0 ;  
                 # 2 0   r e s e t   =   0 ;  
                 f l o o r _ r e q u e s t   =   5 ' b 0 0 0 1 0 ;  
                 # 1 0 0 ;  
                 f l o o r _ r e q u e s t   =   5 ' b 1 0 0 0 0 ;  
                 # 1 0 0 ;  
                 f l o o r _ r e q u e s t   =   5 ' b 0 0 0 1 0 ;  
                 # 1 0 0 ;  
                 f l o o r _ r e q u e s t   =   5 ' b 0 0 0 0 1 ;  
                 # 1 0 0 ;  
                 $ f i n i s h ;  
         e n d  
 e n d m o d u l e 